module pencoder #(
    parameter WIDTH = 6,                     // output width
    parameter DEPTH = (1 << WIDTH) - 1       // number of inputs (32 for WIDTH = 6)
)(
    input [DEPTH-1:0] search_valid_i,
    output reg [WIDTH-1:0] search_index_o
);

always @(*) begin
    casez (search_valid_i)
        32'b????_????_????_????_????_????_????_???1: search_index_o = 6'd0;
        32'b????_????_????_????_????_????_????_??10: search_index_o = 6'd1;
        32'b????_????_????_????_????_????_????_?100: search_index_o = 6'd2;
        32'b????_????_????_????_????_????_????_1000: search_index_o = 6'd3;
        32'b????_????_????_????_????_????_???1_0000: search_index_o = 6'd4;
        32'b????_????_????_????_????_????_??10_0000: search_index_o = 6'd5;
        32'b????_????_????_????_????_????_?100_0000: search_index_o = 6'd6;
        32'b????_????_????_????_????_????_1000_0000: search_index_o = 6'd7;
        32'b????_????_????_????_????_???1_0000_0000: search_index_o = 6'd8;
        32'b????_????_????_????_????_??10_0000_0000: search_index_o = 6'd9;
        32'b????_????_????_????_????_?100_0000_0000: search_index_o = 6'd10;
        32'b????_????_????_????_????_1000_0000_0000: search_index_o = 6'd11;
        32'b????_????_????_????_???1_0000_0000_0000: search_index_o = 6'd12;
        32'b????_????_????_????_??10_0000_0000_0000: search_index_o = 6'd13;
        32'b????_????_????_????_?100_0000_0000_0000: search_index_o = 6'd14;
        32'b????_????_????_????_1000_0000_0000_0000: search_index_o = 6'd15;
        32'b????_????_????_???1_0000_0000_0000_0000: search_index_o = 6'd16;
        32'b????_????_????_??10_0000_0000_0000_0000: search_index_o = 6'd17;
        32'b????_????_????_?100_0000_0000_0000_0000: search_index_o = 6'd18;
        32'b????_????_????_1000_0000_0000_0000_0000: search_index_o = 6'd19;
        32'b????_????_???1_0000_0000_0000_0000_0000: search_index_o = 6'd20;
        32'b????_????_??10_0000_0000_0000_0000_0000: search_index_o = 6'd21;
        32'b????_????_?100_0000_0000_0000_0000_0000: search_index_o = 6'd22;
        32'b????_????_1000_0000_0000_0000_0000_0000: search_index_o = 6'd23;
        32'b????_???1_0000_0000_0000_0000_0000_0000: search_index_o = 6'd24;
        32'b????_??10_0000_0000_0000_0000_0000_0000: search_index_o = 6'd25;
        32'b????_?100_0000_0000_0000_0000_0000_0000: search_index_o = 6'd26;
        32'b????_1000_0000_0000_0000_0000_0000_0000: search_index_o = 6'd27;
        32'b???1_0000_0000_0000_0000_0000_0000_0000: search_index_o = 6'd28;
        32'b??10_0000_0000_0000_0000_0000_0000_0000: search_index_o = 6'd29;
        32'b?100_0000_0000_0000_0000_0000_0000_0000: search_index_o = 6'd30;
        32'b1000_0000_0000_0000_0000_0000_0000_0000: search_index_o = 6'd31;
        default: search_index_o = 6'd32;
    endcase
end

endmodule
